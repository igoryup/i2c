
module unnamed (
	source,
	probe);	

	output	[17:0]	source;
	input	[9:0]	probe;
endmodule
